module coreir_ugt #(parameter width = 1) (input [width-1:0] in0/*verilator public*/, input [width-1:0] in1/*verilator public*/, output out/*verilator public*/);
  assign out = in0 > in1;
endmodule

module coreir_reg #(parameter width = 1, parameter clk_posedge = 1, parameter init = 1) (input clk/*verilator public*/, input [width-1:0] in/*verilator public*/, output [width-1:0] out/*verilator public*/);
  reg [width-1:0] outReg/*verilator public*/=init;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk) begin
    outReg <= in;
  end
  assign out = outReg;
endmodule

module coreir_neg #(parameter width = 1) (input [width-1:0] in/*verilator public*/, output [width-1:0] out/*verilator public*/);
  assign out = -in;
endmodule

module coreir_mux #(parameter width = 1) (input [width-1:0] in0/*verilator public*/, input [width-1:0] in1/*verilator public*/, input sel/*verilator public*/, output [width-1:0] out/*verilator public*/);
  assign out = sel ? in1 : in0;
endmodule

module coreir_const #(parameter width = 1, parameter value = 1) (output [width-1:0] out/*verilator public*/);
  assign out = value;
endmodule

module corebit_and (input in0/*verilator public*/, input in1/*verilator public*/, output out/*verilator public*/);
  assign out = in0 & in1;
endmodule

module top (input CLK/*verilator public*/, output [7:0] O/*verilator public*/, input [7:0] hi/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out;
wire FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$and_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$coreir_const11_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out;
wire FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$and_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$coreir_const11_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out;
wire FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$and_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$coreir_const11_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out;
wire FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$and_inst0_out;
wire [0:0] FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$coreir_const11_inst0_out;
wire [7:0] Map_T_n4_i0_opModule_0_f_in_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0$Module_0_inst0$Abs_Atom_inst0$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out;
wire [7:0] Map_T_n4_i0_opModule_0_f_in_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0$Module_0_inst0$Abs_Atom_inst0$Negate8_inst0$coreir_neg_inst0_out;
wire Map_T_n4_i0_opModule_0_f_in_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0$Module_0_inst0$Abs_Atom_inst0$coreir_ugt8_inst0_out;
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]), .in1(hi[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out[0]), .in1(hi[1]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out[0]), .in1(hi[2]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out[0]), .in1(hi[3]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out[0]), .in1(hi[4]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out[0]), .in1(hi[5]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out[0]), .in1(hi[6]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out[0]), .in1(hi[7]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]), .in1(valid_up), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out));
corebit_and FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$and_inst0(.in0(valid_up), .in1(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$coreir_const11_inst0_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$and_inst0_out));
coreir_const #(.value(1'h1), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$coreir_const11_inst0(.out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$coreir_const11_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]), .in1(Map_T_n4_i0_opModule_0_f_in_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0$Module_0_inst0$Abs_Atom_inst0$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out[0]), .in1(Map_T_n4_i0_opModule_0_f_in_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0$Module_0_inst0$Abs_Atom_inst0$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[1]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out[0]), .in1(Map_T_n4_i0_opModule_0_f_in_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0$Module_0_inst0$Abs_Atom_inst0$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[2]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out[0]), .in1(Map_T_n4_i0_opModule_0_f_in_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0$Module_0_inst0$Abs_Atom_inst0$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[3]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out[0]), .in1(Map_T_n4_i0_opModule_0_f_in_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0$Module_0_inst0$Abs_Atom_inst0$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[4]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out[0]), .in1(Map_T_n4_i0_opModule_0_f_in_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0$Module_0_inst0$Abs_Atom_inst0$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[5]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out[0]), .in1(Map_T_n4_i0_opModule_0_f_in_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0$Module_0_inst0$Abs_Atom_inst0$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[6]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out[0]), .in1(Map_T_n4_i0_opModule_0_f_in_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0$Module_0_inst0$Abs_Atom_inst0$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[7]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]), .in1(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out));
corebit_and FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$and_inst0(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]), .in1(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$coreir_const11_inst0_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$and_inst0_out));
coreir_const #(.value(1'h1), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$coreir_const11_inst0(.out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$coreir_const11_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]), .in1(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out[0]), .in1(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out[0]), .in1(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out[0]), .in1(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out[0]), .in1(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out[0]), .in1(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out[0]), .in1(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out[0]), .in1(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]), .in1(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out));
corebit_and FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$and_inst0(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]), .in1(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$coreir_const11_inst0_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$and_inst0_out));
coreir_const #(.value(1'h1), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$coreir_const11_inst0(.out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$coreir_const11_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]), .in1(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out[0]), .in1(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out[0]), .in1(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out[0]), .in1(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out[0]), .in1(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out[0]), .in1(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out[0]), .in1(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out[0]), .in1(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out));
coreir_mux #(.width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]), .in1(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out), .sel(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$and_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(.clk(CLK), .in(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out));
corebit_and FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$and_inst0(.in0(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]), .in1(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$coreir_const11_inst0_out[0]), .out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$and_inst0_out));
coreir_const #(.value(1'h1), .width(1)) FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$coreir_const11_inst0(.out(FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$coreir_const11_inst0_out));
coreir_mux #(.width(8)) Map_T_n4_i0_opModule_0_f_in_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0$Module_0_inst0$Abs_Atom_inst0$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join(.in0({FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]}), .in1({Map_T_n4_i0_opModule_0_f_in_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0$Module_0_inst0$Abs_Atom_inst0$Negate8_inst0$coreir_neg_inst0_out[7],Map_T_n4_i0_opModule_0_f_in_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0$Module_0_inst0$Abs_Atom_inst0$Negate8_inst0$coreir_neg_inst0_out[6],Map_T_n4_i0_opModule_0_f_in_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0$Module_0_inst0$Abs_Atom_inst0$Negate8_inst0$coreir_neg_inst0_out[5],Map_T_n4_i0_opModule_0_f_in_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0$Module_0_inst0$Abs_Atom_inst0$Negate8_inst0$coreir_neg_inst0_out[4],Map_T_n4_i0_opModule_0_f_in_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0$Module_0_inst0$Abs_Atom_inst0$Negate8_inst0$coreir_neg_inst0_out[3],Map_T_n4_i0_opModule_0_f_in_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0$Module_0_inst0$Abs_Atom_inst0$Negate8_inst0$coreir_neg_inst0_out[2],Map_T_n4_i0_opModule_0_f_in_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0$Module_0_inst0$Abs_Atom_inst0$Negate8_inst0$coreir_neg_inst0_out[1],Map_T_n4_i0_opModule_0_f_in_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0$Module_0_inst0$Abs_Atom_inst0$Negate8_inst0$coreir_neg_inst0_out[0]}), .out(Map_T_n4_i0_opModule_0_f_in_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0$Module_0_inst0$Abs_Atom_inst0$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out), .sel(Map_T_n4_i0_opModule_0_f_in_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0$Module_0_inst0$Abs_Atom_inst0$coreir_ugt8_inst0_out));
coreir_neg #(.width(8)) Map_T_n4_i0_opModule_0_f_in_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0$Module_0_inst0$Abs_Atom_inst0$Negate8_inst0$coreir_neg_inst0(.in({FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]}), .out(Map_T_n4_i0_opModule_0_f_in_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0$Module_0_inst0$Abs_Atom_inst0$Negate8_inst0$coreir_neg_inst0_out));
coreir_ugt #(.width(8)) Map_T_n4_i0_opModule_0_f_in_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0$Module_0_inst0$Abs_Atom_inst0$coreir_ugt8_inst0(.in0({FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]}), .in1(Map_T_n4_i0_opModule_0_f_in_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0$Module_0_inst0$Abs_Atom_inst0$Negate8_inst0$coreir_neg_inst0_out), .out(Map_T_n4_i0_opModule_0_f_in_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0$Module_0_inst0$Abs_Atom_inst0$coreir_ugt8_inst0_out));
assign O = {FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out[0],FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_8_Bit_t_0init_TrueCE_FalseRESET_inst0$Register8CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]};
assign valid_down = FIFO_tTSeq_4_0_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Bitt_0init_TrueCE_FalseRESET_inst0$Register1CE_inst0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0];
endmodule

